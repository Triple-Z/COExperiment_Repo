module mips (clk, rst);
	input clk;
	input rst;

endmodule // mips
