module npc (branch, jump, clk, zero, imm16, ins);
    input branch, jump, clk, zero;
    input      [15:0] imm16;
    output reg [31:0] ins;


endmodule // Next Program Counter;
