library verilog;
use verilog.vl_types.all;
entity pc is
end pc;
