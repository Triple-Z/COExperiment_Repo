module comp();

endmodule // Compare; 