library verilog;
use verilog.vl_types.all;
entity testbench is
end testbench;
