module pc ();

endmodule // Program Counter;
